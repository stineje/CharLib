* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL VSS

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_8 A Y
X0 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X1 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X2 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X3 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X4 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X5 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X6 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X7 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X8 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X9 VDD A a_n8_16 VDD pmos_3p3 w=34 l=6
X10 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X11 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X12 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X13 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X14 VSS A a_n8_16 VSS nmos_3p3 w=17 l=6
X15 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X16 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X17 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
