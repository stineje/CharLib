* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL VSS

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkbuf_16 A Y
X0 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X1 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X2 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X3 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X4 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X5 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X6 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X7 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X8 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X9 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X10 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X11 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X12 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X13 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X14 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X15 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X16 VDD A a_n8_16 VDD pmos_3p3 w=34 l=6
X17 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X18 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
X19 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X20 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X21 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X22 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X23 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X24 VSS a_n8_16 Y VSS nmos_3p3 w=17 l=6
X25 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X26 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X27 VSS A a_n8_16 VSS nmos_3p3 w=17 l=6
X28 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X29 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X30 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X31 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X32 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X33 Y a_n8_16 VSS VSS nmos_3p3 w=17 l=6
C0 VDD Y 2.051450fF
.ends

** hspice subcircuit dictionary
