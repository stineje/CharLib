// Verilog model for OSU350; 
module INVX1(Y,A);
output Y;
input A;
assign Y = !A;
endmodule

